CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 710 30 100 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
36
13 Logic Switch~
5 246 1638 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90098e-315 0
0
13 Logic Switch~
5 195 1423 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90098e-315 0
0
13 Logic Switch~
5 186 1343 0 1 11
0 3
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.90098e-315 0
0
13 Logic Switch~
5 298 1062 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90098e-315 0
0
13 Logic Switch~
5 182 810 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90098e-315 0
0
13 Logic Switch~
5 174 712 0 1 11
0 17
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
5.90098e-315 0
0
13 Logic Switch~
5 114 594 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.90098e-315 0
0
13 Logic Switch~
5 917 488 0 1 11
0 19
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
5.90098e-315 0
0
13 Logic Switch~
5 668 466 0 1 11
0 20
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
5.90098e-315 0
0
13 Logic Switch~
5 472 473 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
5.90098e-315 0
0
13 Logic Switch~
5 242 478 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
5.90098e-315 0
0
13 Logic Switch~
5 186 146 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
5.90098e-315 0
0
14 Logic Display~
6 1060 1308 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
5.90098e-315 0
0
14 Logic Display~
6 845 1293 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
5.90098e-315 0
0
14 Logic Display~
6 664 1287 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
5.90098e-315 0
0
14 Logic Display~
6 449 1282 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.90098e-315 0
0
7 Pulser~
4 121 1746 0 10 12
0 2 29 2 30 0 0 5 5 3
8
0
0 0 4640 0
0
3 V15
-11 -28 10 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5616 0 0
2
5.90098e-315 0
0
5 7474~
219 957 1519 0 6 22
0 3 7 2 9 31 8
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U6B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 6 0
1 U
9323 0 0
2
5.90098e-315 0
0
5 7474~
219 747 1509 0 6 22
0 3 6 2 9 32 7
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U6A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 6 0
1 U
317 0 0
2
5.90098e-315 0
0
5 7474~
219 569 1501 0 6 22
0 3 5 2 9 33 6
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U5B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 5 0
1 U
3108 0 0
2
5.90098e-315 0
0
5 7474~
219 378 1494 0 6 22
0 3 4 2 9 34 5
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U5A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 5 0
1 U
4299 0 0
2
5.90098e-315 0
0
14 Logic Display~
6 1082 761 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.90098e-315 0
0
5 7474~
219 944 953 0 6 22
0 17 15 10 11 35 16
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U4B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 4 0
1 U
7876 0 0
2
5.90098e-315 0
0
5 7474~
219 757 956 0 6 22
0 17 14 10 11 36 15
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U4A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 4 0
1 U
6369 0 0
2
5.90098e-315 0
0
5 7474~
219 539 963 0 6 22
0 17 13 10 11 37 14
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U3B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 3 0
1 U
9172 0 0
2
5.90098e-315 0
0
5 7474~
219 326 957 0 6 22
0 17 12 10 11 38 13
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U3A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 3 0
1 U
7100 0 0
2
5.90098e-315 0
0
7 Pulser~
4 225 1141 0 10 12
0 10 39 10 40 0 0 5 5 3
8
0
0 0 4640 0
0
2 V8
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3820 0 0
2
5.90098e-315 0
0
7 Pulser~
4 60 497 0 10 12
0 18 41 18 42 0 0 5 5 3
8
0
0 0 4640 0
0
2 V7
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7678 0 0
2
5.90098e-315 0
0
14 Logic Display~
6 1104 127 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.90098e-315 0
0
14 Logic Display~
6 888 131 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
5.90098e-315 0
0
14 Logic Display~
6 685 125 0 1 2
10 25
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
5.90098e-315 0
0
14 Logic Display~
6 450 115 0 1 2
10 26
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
5.90098e-315 0
0
5 7474~
219 967 334 0 6 22
0 28 19 18 23 43 27
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 2 0
1 U
8885 0 0
2
5.90098e-315 0
0
5 7474~
219 769 333 0 6 22
0 28 20 18 23 44 24
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 2 0
1 U
3780 0 0
2
5.90098e-315 0
0
5 7474~
219 582 329 0 6 22
0 28 21 18 23 45 25
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 2 1 0
1 U
9265 0 0
2
5.90098e-315 0
0
5 7474~
219 347 318 0 6 22
0 28 22 18 23 46 26
0
0 0 4704 0
4 7474
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
9442 0 0
2
5.90098e-315 0
0
60
3 0 2 0 0 8192 0 19 0 0 3 3
723 1491
693 1491
693 1688
3 0 2 0 0 8192 0 20 0 0 3 3
545 1483
530 1483
530 1688
0 3 2 0 0 4224 0 0 18 20 0 4
131 1688
925 1688
925 1501
933 1501
0 1 3 0 0 4224 0 0 18 5 0 3
747 1440
957 1440
957 1456
0 1 3 0 0 0 0 0 19 6 0 4
569 1405
569 1434
747 1434
747 1446
0 1 3 0 0 0 0 0 20 8 0 3
378 1405
569 1405
569 1438
1 2 4 0 0 4224 0 2 21 0 0 4
207 1423
346 1423
346 1458
354 1458
1 1 3 0 0 0 0 3 21 0 0 3
198 1343
378 1343
378 1431
0 1 5 0 0 4224 0 0 16 10 0 2
449 1458
449 1300
6 2 5 0 0 0 0 21 20 0 0 4
402 1458
537 1458
537 1465
545 1465
0 1 6 0 0 4224 0 0 15 12 0 2
664 1465
664 1305
6 2 6 0 0 0 0 20 19 0 0 4
593 1465
715 1465
715 1473
723 1473
0 1 7 0 0 4224 0 0 14 14 0 2
845 1473
845 1311
6 2 7 0 0 0 0 19 18 0 0 4
771 1473
925 1473
925 1483
933 1483
6 1 8 0 0 8320 0 18 13 0 0 3
981 1483
1060 1483
1060 1326
0 4 9 0 0 4224 0 0 18 17 0 3
747 1554
957 1554
957 1531
0 4 9 0 0 0 0 0 19 18 0 3
569 1560
747 1560
747 1521
0 4 9 0 0 0 0 0 20 19 0 3
378 1566
569 1566
569 1513
1 4 9 0 0 0 0 1 21 0 0 3
258 1638
378 1638
378 1506
0 3 2 0 0 0 0 0 21 21 0 3
131 1723
131 1476
354 1476
1 3 2 0 0 0 0 17 17 0 0 6
97 1737
87 1737
87 1723
159 1723
159 1737
145 1737
3 0 10 0 0 8192 0 25 0 0 24 3
515 945
506 945
506 1089
3 0 10 0 0 8192 0 24 0 0 24 3
733 938
728 938
728 1089
0 3 10 0 0 4224 0 0 23 25 0 4
245 1089
912 1089
912 935
920 935
0 3 10 0 0 0 0 0 26 39 0 3
245 1118
245 939
302 939
0 4 11 0 0 4096 0 0 23 27 0 3
757 973
944 973
944 965
0 4 11 0 0 8320 0 0 24 28 0 4
539 999
539 979
757 979
757 968
0 4 11 0 0 0 0 0 25 29 0 3
326 999
539 999
539 975
1 4 11 0 0 0 0 4 26 0 0 3
310 1062
326 1062
326 969
2 1 12 0 0 8320 0 26 5 0 0 4
302 921
203 921
203 810
194 810
6 2 13 0 0 4224 0 26 25 0 0 4
350 921
507 921
507 927
515 927
6 2 14 0 0 4224 0 25 24 0 0 4
563 927
725 927
725 920
733 920
6 2 15 0 0 4224 0 24 23 0 0 4
781 920
912 920
912 917
920 917
6 1 16 0 0 8320 0 23 22 0 0 3
968 917
1082 917
1082 779
0 1 17 0 0 4096 0 0 23 36 0 3
757 861
944 861
944 890
0 1 17 0 0 4224 0 0 24 37 0 3
539 851
757 851
757 893
0 1 17 0 0 0 0 0 25 38 0 3
326 844
539 844
539 900
1 1 17 0 0 0 0 6 26 0 0 3
186 712
326 712
326 894
1 3 10 0 0 0 0 27 27 0 0 6
201 1132
191 1132
191 1118
263 1118
263 1132
249 1132
0 3 18 0 0 4096 0 0 35 42 0 3
514 436
514 311
558 311
0 3 18 0 0 0 0 0 34 42 0 3
703 436
703 315
745 315
0 3 18 0 0 4224 0 0 33 43 0 4
63 436
930 436
930 316
943 316
0 3 18 0 0 0 0 0 36 52 0 3
63 474
63 300
323 300
1 2 19 0 0 8320 0 8 33 0 0 4
929 488
935 488
935 298
943 298
1 2 20 0 0 8320 0 9 34 0 0 4
680 466
737 466
737 297
745 297
1 2 21 0 0 8320 0 10 35 0 0 4
484 473
550 473
550 293
558 293
1 2 22 0 0 8320 0 11 36 0 0 4
254 478
315 478
315 282
323 282
1 0 23 0 0 8320 0 7 0 0 55 3
126 594
369 594
369 349
6 1 24 0 0 8320 0 34 30 0 0 3
793 297
888 297
888 149
6 1 25 0 0 8320 0 35 31 0 0 3
606 293
685 293
685 143
6 1 26 0 0 8320 0 36 32 0 0 3
371 282
450 282
450 133
1 3 18 0 0 0 0 28 28 0 0 6
36 488
26 488
26 474
98 474
98 488
84 488
0 4 23 0 0 0 0 0 33 54 0 4
768 353
768 359
967 359
967 346
0 4 23 0 0 0 0 0 34 55 0 4
580 349
580 353
769 353
769 345
4 4 23 0 0 0 0 36 35 0 0 4
347 330
347 349
582 349
582 341
6 1 27 0 0 8320 0 33 29 0 0 3
991 298
1104 298
1104 145
0 1 28 0 0 4096 0 0 33 58 0 3
769 195
967 195
967 271
0 1 28 0 0 0 0 0 34 59 0 3
582 186
769 186
769 270
0 1 28 0 0 4224 0 0 35 60 0 3
347 179
582 179
582 266
1 1 28 0 0 0 0 12 36 0 0 3
198 146
347 146
347 255
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
522 1156 607 1180
532 1164 596 1180
8 FIG:SISO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
426 621 511 645
436 629 500 645
8 Fig:PIPO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
454 1798 539 1822
464 1806 528 1822
8 Fig:SIPO
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
